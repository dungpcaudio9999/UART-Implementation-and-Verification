`timescale 1ns/1ps

module tb_uart_core;

    // =========================================================================
    // 1. SIGNALS & CONSTANTS
    // =========================================================================
    // Clock & Reset
    reg clk;
    reg rst_n;
    
    // Configuration
    reg [15:0] i_divisor;
    reg [1:0]  i_num_bit_data;
    reg        i_parity_en;
    reg        i_parity_type; // 0: Even, 1: Odd

    // CPU Interface
    reg [7:0]  i_cpu_txd;
    reg        i_tx_wr;
    wire       o_tx_full;
    wire [7:0] o_cpu_rxd;
    reg        i_rx_rd;
    wire       o_rx_empty;
    wire       o_parity_err;

    // Physical Interface
    wire       o_pedev_txd;
    reg        i_pedev_rxd;
    reg        i_cts_n;
    wire       o_rts_n;

    // Testbench Control Signals
    reg        loopback_en; // 1: Internal Loopback, 0: External Stimulus
    reg        stim_rxd;    // Generated by TB task

    // capture parity error
    reg parity_err_latched;

    // Constants for 50MHz Clock
    localparam CLK_PERIOD = 20; 
    
    // =========================================================================
    // 2. DUT INSTANTIATION [cite: 30]
    // =========================================================================
    uart_core dut (
        .clk            (clk),
        .rst_n          (rst_n),
        .i_divisor      (i_divisor),
        .i_num_bit_data (i_num_bit_data),
        .i_parity_en    (i_parity_en),
        .i_parity_type  (i_parity_type),
        .i_cpu_txd      (i_cpu_txd),
        .i_tx_wr        (i_tx_wr),
        .o_tx_full      (o_tx_full),
        .o_cpu_rxd      (o_cpu_rxd),
        .i_rx_rd        (i_rx_rd),
        .o_rx_empty     (o_rx_empty),
        .o_parity_err   (o_parity_err),
        .o_pedev_txd    (o_pedev_txd),
        .i_pedev_rxd    (i_pedev_rxd),
        .i_cts_n        (i_cts_n),
        .o_rts_n        (o_rts_n)
    );

    // Loopback Mux Logic
    always @(loopback_en or o_pedev_txd or stim_rxd) begin
        if (loopback_en)
            i_pedev_rxd = o_pedev_txd;
        else
            i_pedev_rxd = stim_rxd;
    end

    // Logic: capture o_parity_err 
    always @(posedge clk) begin
        if (o_parity_err) 
            parity_err_latched <= 1'b1;
    end

    // Clock Generation
    initial begin
        clk = 0;
        forever #(CLK_PERIOD/2) clk = ~clk;
    end

    // =========================================================================
    // 3. TASKS
    // =========================================================================
    
    // Task: Reset System
    task apply_reset();
        begin
            rst_n = 0;
            i_tx_wr = 0;
            i_rx_rd = 0;
            i_cts_n = 0; // Clear to send active (Low)
            loopback_en = 0;
            stim_rxd = 1;
            i_divisor = 325; // Default 9600
            i_num_bit_data = 2'b11; // 8 bits
            i_parity_en = 0;
            i_parity_type = 0;
            repeat(5) @(posedge clk);
            rst_n = 1;
            @(posedge clk);
        end
    endtask

    // Task: CPU Write to TX FIFO
    task cpu_write(input [7:0] data);
        begin
            @(posedge clk);
            while(o_tx_full) @(posedge clk); // Wait if full (optional flow control)
            i_cpu_txd = data;
            i_tx_wr = 1;
            @(posedge clk);
            i_tx_wr = 0;
        end
    endtask

    // Task: CPU Read from RX FIFO
    task cpu_read(output [7:0] data);
    begin
        @(posedge clk);
        // Wait for data
        while(o_rx_empty) @(posedge clk);
        i_rx_rd = 1;
        data = o_cpu_rxd; // Capture data
        @(posedge clk); // Allow FIFO to update output

        i_rx_rd = 0;
    end
    endtask

    // Task: Simulate External UART Device sending to DUT
    task drive_rx_serial(
        input [7:0] data,
        input       inject_parity_err
    );
        integer i;
        reg parity_bit;
        integer bit_width;
        integer bit_ticks;
        begin
            // Calculate bit timing
            bit_ticks = i_divisor * 16;     // RX need 16 tick
            
            // Calculate effective data width
            case(i_num_bit_data)
                2'b00: bit_width = 5;
                2'b01: bit_width = 6;
                2'b10: bit_width = 7;
                2'b11: bit_width = 8;
            endcase

            // Calculate Parity
            parity_bit = 0;
            case(i_num_bit_data)
                2'b00: parity_bit = ^data[4:0];
                2'b01: parity_bit = ^data[5:0];
                2'b10: parity_bit = ^data[6:0];
                2'b11: parity_bit = ^data[7:0];
            endcase
            
            if(i_parity_type) parity_bit = ~parity_bit; // Odd parity
            if(inject_parity_err) parity_bit = ~parity_bit; // Force Error

            // --- Start Transmission ---
            // 1. Start Bit (Low)
            stim_rxd = 0;
            repeat(bit_ticks) @(posedge clk);

            // 2. Data Bits (LSB first)
            for(i=0; i<bit_width; i=i+1) begin
                stim_rxd = data[i];
                repeat(bit_ticks) @(posedge clk);
            end

            // 3. Parity Bit (Optional)
            if(i_parity_en) begin
                stim_rxd = parity_bit;
                repeat(bit_ticks) @(posedge clk);
            end

            // 4. Stop Bit (High)
            stim_rxd = 1;
            repeat(bit_ticks) @(posedge clk);
        end
    endtask

    // Helper: Wait for n baud periods
    task wait_baud_periods(input integer n);
        repeat(n * 16 * i_divisor) @(posedge clk);
    endtask

    // =========================================================================
    // 4. MAIN TEST SEQUENCE
    // =========================================================================
    reg [7:0] read_val;
    integer k;

    initial begin
        // Setup waveforms
        $dumpfile("uart_dump.vcd");
        $dumpvars(0, tb_uart_core);

        $display("----------------------------------------------------------------");
        $display("STARTING UART VERIFICATION");
        $display("----------------------------------------------------------------");

        apply_reset();

        // ---------------------------------------------------------------------
        // CORE_01: Sanity - Internal Loopback
        // ---------------------------------------------------------------------
        $display("[CORE_01] Sanity: Internal Loopback (9600, 8N1)");
        i_divisor = 325; // 9600
        i_num_bit_data = 2'b11; // 8 bit
        i_parity_en = 0;
        loopback_en = 1;
        
        cpu_write(8'hA5);
        $display("[DEBUG] rx empty value: %b", o_rx_empty);
        $display("[DEBUG] Read value: %0h", read_val);
        
        // Wait enough time for TX -> RX
        wait_baud_periods(12);
        $display("[DEBUG] Read value: %0h", read_val);
        $display("[DEBUG] rx empty value: %b", o_rx_empty); 
        
        if(o_rx_empty == 0) begin
            $display("[DEBUG] Read value: %0h", read_val);
            cpu_read(read_val);
            $display("[DEBUG] Read value: %0h", read_val);
            if(read_val == 8'hA5) $display("  -> PASSED: Received 0xA5");
            else $error("  -> FAILED: Expected 0xA5, got 0x%h", read_val);
        end else begin
            $error("  -> FAILED: RX FIFO Empty (Timeout)");
        end

        // ---------------------------------------------------------------------
        // CORE_02: TX Path - FIFO TX Full Flag
        // ---------------------------------------------------------------------
        $display("\n[CORE_02] TX Path: TX FIFO Full Flag");
        loopback_en = 0; // Disconnect RX to verify TX only
        // To test FULL, we need to fill faster than TX can drain.
        // Or block CTS. Let's block CTS to keep data in FIFO.
        i_cts_n = 1; 
        
        // FIFO Depth is 16. Write 16 bytes.
        for(k=0; k<16; k=k+1) begin
            cpu_write(8'h00 + k);
        end
        
        // Check Full Flag
        @(posedge clk);
        if(o_tx_full == 1'b1) $display("  -> PASSED: FIFO Full Flag Asserted after 16 bytes");
        else $error("  -> FAILED: FIFO Full Flag not asserted (Status: %b)", o_tx_full);

        i_cts_n = 0; // Release CTS
        wait_baud_periods(20); // Let it drain a bit

        // ---------------------------------------------------------------------
        // CORE_03: TX Path - FIFO TX Empty Flag
        // ---------------------------------------------------------------------
        $display("\n[CORE_03] TX Path: FIFO TX Empty Flag");
        // Wait until all data drains
        wait_baud_periods(16 * 11); 
        
        // Use hierarchical reference to check internal FIFO empty signal 
        // because uart_core doesn't expose o_tx_empty to CPU, only o_tx_full.
        if(dut.u_tx_fifo.o_empty == 1'b1) 
            $display("  -> PASSED: Internal TX FIFO Empty Flag Asserted");
        else 
            $error("  -> FAILED: Internal TX FIFO not empty");

        // ---------------------------------------------------------------------
        // CORE_04: RX Path - Receive & Read
        // ---------------------------------------------------------------------
        $display("\n[CORE_04] RX Path: Receive & Read 0x55");
        loopback_en = 0;
        i_num_bit_data = 2'b11; // 8N1
        i_parity_en = 0;
        
        drive_rx_serial(8'h55, 0); // Send 0x55
        $display("[DEBUG] Read value: %0h", read_val);
        $display("[DEBUG] rx empty value: %b", o_rx_empty); 
        
        @(posedge clk);
        if(o_rx_empty == 0) begin
            cpu_read(read_val);
            if(read_val == 8'h55) $display("  -> PASSED: Read 0x55 correctly");
            else $error("  -> FAILED: Expected 0x55, got 0x%h", read_val);
        end else $error("  -> FAILED: RX FIFO Empty");

        // ---------------------------------------------------------------------
        // CORE_05: RX Path - Parity Check (Good)
        // ---------------------------------------------------------------------
        $display("\n[CORE_05] RX Path: Parity Check (Good) - 8-Even-1");
        i_num_bit_data = 2'b11; 
        i_parity_en = 1;
        i_parity_type = 0; // Even
        
        // Send 0x03 (Bin: 00000011). Even parity -> Parity Bit = 0.
        // drive_rx_serial calculates this automatically.
        drive_rx_serial(8'h03, 0); 
        
        @(posedge clk);
        cpu_read(read_val); // Clear FIFO
        if(o_parity_err === 0 && read_val === 8'h03) 
            $display("  -> PASSED: Data 0x03 received, No Parity Error");
        else 
            $error("  -> FAILED: Err=%b, Data=0x%h", o_parity_err, read_val);

        // ---------------------------------------------------------------------
        // CORE_06: RX Path - Parity Check (Bad)
        // ---------------------------------------------------------------------
        $display("\n[CORE_06] RX Path: Parity Check (Bad) - 8-Even-1");
        i_num_bit_data = 2'b11;
        i_parity_en = 1;     // Enable Parity
        i_parity_type = 0;   // Even

        // delete parity flag before test
        parity_err_latched = 0;

        // Send 0x03 but force error injection
        drive_rx_serial(8'h03, 1);
        $display("[DEBUG] parity error: %b", parity_err_latched); 
        
        @(posedge clk);
        // Note: o_parity_err updates immediately upon RX Done
        $display("[DEBUG] parity error: %b", parity_err_latched);
        if(parity_err_latched == 1) 
            $display("  -> PASSED: Parity Error Flag detected");
        else 
            $error("  -> FAILED: Parity Error Flag NOT detected");
        
        // Read to clear for next test
        if(!o_rx_empty) cpu_read(read_val);

        // ---------------------------------------------------------------------
        // CORE_07: Config - Baud Rate Change (19200)
        // ---------------------------------------------------------------------
        $display("\n[CORE_07] Config: Baud Rate Change to 19200");
        loopback_en = 1;
        i_parity_en = 0;
        i_divisor = 162; // 19200bps @ 50MHz
        
        cpu_write(8'hCC);
        
        // Wait shorter time (since faster baud)
        wait_baud_periods(12);
        
        if(!o_rx_empty) begin
            cpu_read(read_val);
            if(read_val === 8'hCC) $display("  -> PASSED: Loopback 0xCC at 19200bps");
            else $error("  -> FAILED: Data mismatch 0x%h", read_val);
        end else $error("  -> FAILED: No data received");

        // ---------------------------------------------------------------------
        // CORE_08: Config - Data Width (5-bit)
        // ---------------------------------------------------------------------
        $display("\n[CORE_08] Config: Data Width 5-bit");
        i_divisor = 325; // Back to 9600
        i_num_bit_data = 2'b00; // 5 bits
        
        cpu_write(8'h1F); // 0001 1111 (All 5 bits high)
        wait_baud_periods(12);
        
        if(!o_rx_empty) begin
            cpu_read(read_val);
            // Expect upper 3 bits to be 0
            if(read_val === 8'h1F) $display("  -> PASSED: Received 0x1F in 5-bit mode");
            else $error("  -> FAILED: Expected 0x1F, got 0x%h", read_val);
        end

        // ---------------------------------------------------------------------
        // CORE_09: Flow Ctrl - RTS Trigger
        // ---------------------------------------------------------------------
        $display("\n[CORE_09] Flow Ctrl: RTS Trigger");
        loopback_en = 0;
        i_num_bit_data = 2'b11; // 8 bit
        
        // Reset RX FIFO to be empty first
        apply_reset(); 
        
        // Inject 14 bytes rapidly without reading
        $display("  -> Injecting 14 bytes...");
        for(k=0; k<14; k=k+1) begin
            drive_rx_serial(8'hA0 + k, 0);
        end
        
        // Check RTS. Code says o_rts_n = rx_fifo_almost_full
        // If Almost Full (>=14), o_rts_n should be 1.
        @(posedge clk);
        if(o_rts_n === 1'b1) $display("  -> PASSED: RTS asserted (High) after 14 bytes");
        else $error("  -> FAILED: RTS is %b (Expected 1)", o_rts_n);

        // ---------------------------------------------------------------------
        // CORE_10: Flow Ctrl - CTS Blocking
        // ---------------------------------------------------------------------
        $display("\n[CORE_10] Flow Ctrl: CTS Blocking");
        // Reset to clear state
        apply_reset();
        
        i_cts_n = 1; // Assert CTS (Active High blocking as per logic observed in CORE_02/Code)
                     // Wait, code maps .i_cts_n(i_cts_n).
                     // Code in uart_tx: if(i_tx_start && !i_cts_n)
                     // So !i_cts_n must be TRUE to start. i_cts_n must be 0 to start.
                     // If i_cts_n = 1, it blocks.
        
        cpu_write(8'hAA);
        
        // Wait 1 baud period. TX line should remain IDLE (1).
        wait_baud_periods(1);
        
        if(o_pedev_txd === 1'b1) 
            $display("  -> PASSED: TX Line held IDLE while CTS is High");
        else 
            $error("  -> FAILED: TX Line toggled low despite CTS blocking");

        // Release CTS and see if it sends
        i_cts_n = 0;
        @(posedge clk);
        wait_baud_periods(1);
        if(o_pedev_txd === 1'b0) // Start bit
            $display("  -> PASSED: Transmission started after CTS released");
        
        $display("----------------------------------------------------------------");
        $display("TEST COMPLETED");
        $display("----------------------------------------------------------------");
        $finish;
    end

endmodule